module magy

pub fn hello() {
	cat('dd')
}
