module magy
